module constant_value_generator #(parameter W=32, val=7) (output [W-1:0] out);

assign out= val;

endmodule